
--Updated on March 26th, 2014 
--Changes
--------------------------------------------- 
--Added additional input port clock
--Removed byte-wise reading and writing
----------------------------------------------
--Updated on March 29th, 2014
--Changes
--------------------------------------------- 
--ignoring the 2 LSBs of address
--incresed memory depth to avoid out of bounds for
----address
----------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all;

entity datamem is
    Port ( clock      : in std_logic;
	       address, ext_addr    : in  STD_LOGIC_VECTOR (31 downto 0);
           write_data : in  STD_LOGIC_VECTOR (31 downto 0);
           MemWrite   : in  STD_LOGIC;
           MemRead    : in  STD_LOGIC;
           Read_data, ext_read  : out  STD_LOGIC_VECTOR (31 downto 0));
end datamem;

architecture Behavioral of datamem is
type datamem1 is array (0 to 19199) of std_logic_vector (31 downto 0);
--signal a1,a2,a3,a4:std_logic_vector(5 downto 0);
signal data_out:std_logic_vector(31 downto 0);
signal RAM: datamem1:=(
	x"00000000", -- frame buffer
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"ffffffff", -- image
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fff00001",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ff800000",
	x"3fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fc000000",
	x"01ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"f0000000",
	x"007fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"c0000000",
	x"001fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"80000000",
	x"0007ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"00000000",
	x"0000ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffffe",
	x"00000000",
	x"00007fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffffc",
	x"00000000",
	x"00001fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff8",
	x"00000000",
	x"00000fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff0",
	x"00000000",
	x"000007ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff0",
	x"0000fff0",
	x"000001ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff0",
	x"0007ffff",
	x"800000ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff0",
	x"001fffff",
	x"e000007f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff0",
	x"003fffff",
	x"f800001f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff0",
	x"003fffff",
	x"fe00000f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff0",
	x"003fffff",
	x"ff800007",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff0",
	x"003fffff",
	x"ffc00003",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff0",
	x"001fffff",
	x"ffe00003",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff0",
	x"000fffff",
	x"fff80001",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff0",
	x"000fffff",
	x"fffc0000",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff8",
	x"0007ffff",
	x"fffe0000",
	x"7fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff8",
	x"0003ffff",
	x"ffff0000",
	x"3fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffffc",
	x"0001ffff",
	x"ffff8000",
	x"1fffffff",
	x"fffffff8",
	x"003fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffffe",
	x"0001ffff",
	x"ffffc000",
	x"0fffffff",
	x"fffffe00",
	x"0003ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffffe",
	x"0000ffff",
	x"ffffe000",
	x"07ffffff",
	x"fff80000",
	x"00001fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"00007fff",
	x"fffff000",
	x"07ffffff",
	x"ffc00000",
	x"000007ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"80003fff",
	x"fffff800",
	x"03ffffff",
	x"f0000000",
	x"000003ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"80001fff",
	x"fffffc00",
	x"01ffffff",
	x"80000000",
	x"000000ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"c00007ff",
	x"fffffe00",
	x"00fffffc",
	x"00000000",
	x"000000ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"e00003ff",
	x"ffffff00",
	x"00ffffc0",
	x"00000000",
	x"0000007f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"f00001ff",
	x"ffffff00",
	x"007fff00",
	x"00000000",
	x"0000003f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"f80000ff",
	x"ffffff80",
	x"003fe000",
	x"00000000",
	x"0000003f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fc00007f",
	x"ffffffc0",
	x"001f8000",
	x"00000000",
	x"0000003f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fe00001f",
	x"ffffffe0",
	x"00000000",
	x"00000000",
	x"0000003f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ff00000f",
	x"ffffffe0",
	x"00000000",
	x"00000fff",
	x"ff00001f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffc00007",
	x"fffffff0",
	x"00000000",
	x"00007fff",
	x"ff80001f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffe00003",
	x"fffffff8",
	x"00000000",
	x"000fffff",
	x"ffc0001f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffe00001",
	x"fffffffc",
	x"00000000",
	x"007fffff",
	x"ffe0001f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffe00000",
	x"fffffffc",
	x"00000000",
	x"0fffffff",
	x"ffe0001f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ff800000",
	x"7ffffffc",
	x"00000000",
	x"7fffffff",
	x"ffe0001f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fc000000",
	x"3ffffffc",
	x"00000003",
	x"ffffffff",
	x"ffe0001f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff8",
	x"00000000",
	x"03fffffe",
	x"0000003f",
	x"ffffffff",
	x"ffe0003f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffff80",
	x"00000000",
	x"01ffffff",
	x"000001ff",
	x"ffffffff",
	x"ffc0003f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff800",
	x"00000000",
	x"007fffff",
	x"800007ff",
	x"ffffffff",
	x"ff80007f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff8000",
	x"00000000",
	x"003fffff",
	x"c0001fff",
	x"ffffffff",
	x"fe0000ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffc0000",
	x"00000000",
	x"001fffff",
	x"e0003fff",
	x"ffffffff",
	x"fc0000ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ff000000",
	x"00000000",
	x"001fffff",
	x"f800ffff",
	x"ffffffff",
	x"f00000ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fc000000",
	x"00000000",
	x"001fffff",
	x"fe01ffff",
	x"ffffffff",
	x"c00001ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"80000000",
	x"00000000",
	x"003fffff",
	x"ffcfffff",
	x"ffffffff",
	x"000003ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"00000000",
	x"00000000",
	x"007fffff",
	x"ffffffff",
	x"fffffffc",
	x"000007ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff0",
	x"00000000",
	x"00000000",
	x"00ffffff",
	x"ffffffff",
	x"fffffff0",
	x"00000fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffc0",
	x"00000000",
	x"07ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffff80",
	x"00001fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffff00",
	x"00000000",
	x"3fffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffe00",
	x"00007fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff800",
	x"0000001f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff800",
	x"0001ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffe000",
	x"000000ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffc000",
	x"0003ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff0000",
	x"00000fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff0000",
	x"000fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fff80000",
	x"0001ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffc0000",
	x"001fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fff00000",
	x"0007ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fff80000",
	x"007fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ff800000",
	x"00ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fff00000",
	x"007fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fe000000",
	x"07ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fff00000",
	x"007fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"f8000000",
	x"3fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fff00000",
	x"001fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"f0000000",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fff00000",
	x"0003ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"e0000001",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fff80000",
	x"0000ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"80000007",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffc0000",
	x"00000fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"0000003f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffe0000",
	x"000003ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffffc",
	x"000000ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff0000",
	x"0000000f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff8",
	x"000003ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffe000",
	x"00000001",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffe0",
	x"00000fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff800",
	x"00000000",
	x"07ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffff80",
	x"0000ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffc0",
	x"00000000",
	x"01ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffe00",
	x"003fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"00000000",
	x"001fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff800",
	x"0fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"f8000000",
	x"0003ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff000",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ff000000",
	x"0000ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffc007",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffc00000",
	x"00003fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff803f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fff80000",
	x"00000fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffe00ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff0000",
	x"000003ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffc03ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff000",
	x"000001ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fff007ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffff00",
	x"0000007f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffc00fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffffc",
	x"0000003f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ff001fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"8000001f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fe007fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"f0000007",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"f800ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fe000003",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"f001ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ff800000",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"e001ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffe00000",
	x"7fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"8003ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffc0000",
	x"3fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"0007ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff0000",
	x"1fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffffe",
	x"0007ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff8000",
	x"0fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffffc",
	x"000fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffc000",
	x"07ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff0",
	x"000fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffe000",
	x"03ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffe0",
	x"000fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff800",
	x"01ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffc0",
	x"001fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff800",
	x"007fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffff00",
	x"001fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffc00",
	x"003fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffe00",
	x"003fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffff00",
	x"001fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffc00",
	x"007fffff",
	x"ffffffff",
	x"fffffffe",
	x"000007ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffff80",
	x"0007ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff000",
	x"00ffffff",
	x"ffffffff",
	x"fffffff0",
	x"000000ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffc0",
	x"0003ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffe000",
	x"03ffffff",
	x"ffffffff",
	x"ffffffe0",
	x"0000007f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffe0",
	x"0001ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff8000",
	x"07ffffff",
	x"ffffffff",
	x"ffffffc0",
	x"0000003f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff0",
	x"0000ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff0000",
	x"0fffffff",
	x"ffffffff",
	x"ffffff80",
	x"0000001f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffffc",
	x"00003fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffe0000",
	x"3fffffff",
	x"ffffffff",
	x"ffffff80",
	x"0000001f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffffe",
	x"00001fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffc0000",
	x"7fffffff",
	x"ffffffff",
	x"ffffff00",
	x"0000001f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"00000fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fff00000",
	x"ffffffff",
	x"ffffffff",
	x"ffffff00",
	x"0000003f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"c00003ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffe00003",
	x"ffffffff",
	x"ffffffff",
	x"ffffff00",
	x"0000003f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"e00001ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffc00007",
	x"ffffffff",
	x"ffffffff",
	x"ffffff00",
	x"000000ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"f00000ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ff00000f",
	x"ffffffff",
	x"ffffffff",
	x"ffffff80",
	x"000003ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fc00007f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fe00001f",
	x"ffffffff",
	x"ffffffff",
	x"ffffff80",
	x"00000fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fe00001f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"f800007f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffc0",
	x"0003ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ff00000f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"f00000ff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff0",
	x"003fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ff800007",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"c00001ff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff8",
	x"00ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffe00001",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"800007ff",
	x"ffffffff",
	x"ffffffff",
	x"fffffffe",
	x"0fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fff00000",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"00000fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fff80000",
	x"7fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffffc",
	x"00001fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffe0000",
	x"1fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff8",
	x"00007fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff0000",
	x"0fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffe0",
	x"0001ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffc000",
	x"07ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffff80",
	x"0003ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffe000",
	x"03ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffe00",
	x"0007ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff000",
	x"00ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff800",
	x"000fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff800",
	x"00ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff000",
	x"003fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffc00",
	x"003fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffc000",
	x"007fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffff00",
	x"003fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff8000",
	x"00ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffff80",
	x"001fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff0000",
	x"03ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffc0",
	x"000fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffc0000",
	x"07ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffe0",
	x"0007ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fff80000",
	x"1fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff0",
	x"0001ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fff00000",
	x"3fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff8",
	x"0000ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffe00000",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffffc",
	x"00007fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ff800001",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffffe",
	x"00003fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ff000007",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"c3ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"00001fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fe00000f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffffc",
	x"007fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"80000fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fc00007f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffe0",
	x"001fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"e00007ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"f00000ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffff80",
	x"000fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"f00007ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"e00003ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffe00",
	x"0007ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"f80003ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"e00007ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffe000",
	x"0007ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fc0001ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"c0000fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff0000",
	x"0007ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fc0000ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"80001fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fff00000",
	x"000fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fe0000ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"00003fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ff800000",
	x"001fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ff00007f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffffe",
	x"00003fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"f8000000",
	x"007fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ff80003f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffffe",
	x"0000ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"c0000000",
	x"03ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffc0001f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffffc",
	x"0001ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff8",
	x"00000000",
	x"7fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffe0001f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff8",
	x"0003ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffe0",
	x"00000003",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffe0000f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff8",
	x"0007ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff800",
	x"0000003f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fff0000f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff8",
	x"000fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffe000",
	x"000001ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fff80003",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff8",
	x"000fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffc0000",
	x"00003fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffc0003",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff0",
	x"001fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffe00000",
	x"0001ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffc0003",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff0",
	x"001fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fe000000",
	x"003fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffe0001",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff0",
	x"003fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"e0000000",
	x"00ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff0000",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff0",
	x"003fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"80000000",
	x"3fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff8000",
	x"7fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff0",
	x"003fffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff8",
	x"00000000",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff8000",
	x"7fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff0",
	x"001fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffc0",
	x"0000000f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffc000",
	x"3fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff0",
	x"000fffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff000",
	x"0000003f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffc000",
	x"3fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff0",
	x"000fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff8000",
	x"000003ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffe000",
	x"1fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff8",
	x"0007ffff",
	x"ffffffff",
	x"ffffffff",
	x"ff800000",
	x"000007ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff000",
	x"0fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff8",
	x"0003ffff",
	x"ffffffff",
	x"ffffffff",
	x"fc000000",
	x"00001fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff000",
	x"0fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff8",
	x"0001ffff",
	x"ffffffff",
	x"fffffff0",
	x"00000000",
	x"00001fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff000",
	x"0fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff8",
	x"00007fff",
	x"ffffffff",
	x"ffffffc0",
	x"00000000",
	x"00001fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff800",
	x"07ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffffc",
	x"000007ff",
	x"ffffffff",
	x"fffe0000",
	x"00000000",
	x"00001fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff800",
	x"07ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffffe",
	x"0000007f",
	x"ffffffff",
	x"fff00000",
	x"00000000",
	x"00000fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffc00",
	x"03ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"80000000",
	x"0fffffff",
	x"80000000",
	x"00000000",
	x"00000fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffe00",
	x"01ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"c0000000",
	x"000fff80",
	x"00000000",
	x"00000000",
	x"000007ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffe00",
	x"01ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"e0000000",
	x"00000000",
	x"00000000",
	x"0000003f",
	x"000007ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffff00",
	x"01ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"f8000000",
	x"00000000",
	x"00000000",
	x"000007ff",
	x"000007ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffff00",
	x"00ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fc000000",
	x"00000000",
	x"00000000",
	x"00003fff",
	x"800003ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffff80",
	x"007fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ff000000",
	x"00000000",
	x"00000000",
	x"0007ffff",
	x"800003ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffc0",
	x"007fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ff800000",
	x"00000000",
	x"00000000",
	x"007fffff",
	x"c00003ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffc0",
	x"007fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffe00000",
	x"00000000",
	x"00000000",
	x"03ffffff",
	x"c00003ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffc0",
	x"003fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fff80000",
	x"00000000",
	x"0000003f",
	x"ffffffff",
	x"e00003ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffe0",
	x"003fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff0000",
	x"00000000",
	x"000001ff",
	x"ffffffff",
	x"e00007ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffe0",
	x"001fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffff80",
	x"00000000",
	x"0007ffff",
	x"ffffffff",
	x"e00007ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff0",
	x"000fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffffc",
	x"00000000",
	x"007fffff",
	x"ffffffff",
	x"e00007ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff8",
	x"000fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ff80000f",
	x"ffffffff",
	x"ffffffff",
	x"e0000fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff8",
	x"0007ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"e0001fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff8",
	x"0003ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"e0001fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffffc",
	x"0001ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"f0001fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffffe",
	x"00007fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"f8000fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffffe",
	x"00001fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"f8000fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"00000fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"f80007ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"000007ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fc0007ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"000007ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fc0007ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"800007ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fc0003ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"c00007ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fe0003ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"c00007ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ff0001ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"e00007ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ff0001ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"e00007ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ff0000ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"f00007ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ff8000ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"f80007ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ff8000ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"f80007ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ff80007f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"f80003ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffc0007f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fc0003ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffe0003f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fc0001ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffe0003f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fe0000ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffe0001f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ff0000ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fff0001f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ff0000ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fff0001f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ff80007f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fff8000f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffc0003f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fff8000f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffc0003f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffc0007",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffe0001f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffc0003",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fff0001f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffc0003",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fff0000f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffc0003",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fff80007",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffe0003",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fff80003",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffe0001",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffc0003",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff0001",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffc0003",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff8000",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffc0003",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff8000",
	x"7fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffc0003",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff8000",
	x"7fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffc0003",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff8000",
	x"7fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffc0003",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffc000",
	x"7fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffc0003",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffc000",
	x"7fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffc0003",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffc000",
	x"7fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffc0003",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffe000",
	x"7fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffc0003",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffe000",
	x"7fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffc0003",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff000",
	x"3fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffc0003",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff000",
	x"1fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffc0003",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff000",
	x"1fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffc0003",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff000",
	x"0fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffc0003",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff000",
	x"0fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffc0003",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff000",
	x"0fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffc0003",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff000",
	x"0fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffe0003",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff000",
	x"0fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffe0003",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff800",
	x"0fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff0003",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff800",
	x"0fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff0003",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff800",
	x"0fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff0003",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff800",
	x"0fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff8003",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff800",
	x"0fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff8003",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff800",
	x"0fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff8001",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff800",
	x"0fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff8001",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff800",
	x"0fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff8001",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff000",
	x"0fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff8001",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffc000",
	x"0fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff8000",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"c0000000",
	x"0fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff8000",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffffc",
	x"00000000",
	x"0fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff8000",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffe0",
	x"00000000",
	x"0fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff8000",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffe00",
	x"00000000",
	x"0fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff8000",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffe0",
	x"00000000",
	x"00000000",
	x"0fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff8000",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffc00",
	x"00000000",
	x"00000000",
	x"1fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff8000",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff8000",
	x"00000000",
	x"00000000",
	x"3fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff8000",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffe00000",
	x"00000000",
	x"00000000",
	x"7fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff8000",
	x"7fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ff800000",
	x"00000000",
	x"00000001",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffc000",
	x"7fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ff000000",
	x"00000000",
	x"00000003",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffc000",
	x"7fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fe000000",
	x"00000000",
	x"0000003f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffe000",
	x"7fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"f8000000",
	x"00000000",
	x"000007ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffe000",
	x"3fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"f0000000",
	x"00000000",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffe000",
	x"1fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"f0000000",
	x"00000003",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff000",
	x"1fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"e0000000",
	x"000000ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff000",
	x"0fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"c0000000",
	x"000007ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff000",
	x"0fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"c00001ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff800",
	x"0fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"c0000fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffc00",
	x"0fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"c0001fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffc00",
	x"07ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"c0003fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffc00",
	x"03ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"c0007fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffc00",
	x"03ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"c0007fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffc00",
	x"03ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"c0007fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffc00",
	x"03ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"c0007fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffc00",
	x"03ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"c0003fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffe00",
	x"03ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"c0001fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffe00",
	x"03ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"c00003ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffc00",
	x"03ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"c000000f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffc00",
	x"03ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"e0000000",
	x"0007ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffc00",
	x"03ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"f0000000",
	x"0000ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffc00",
	x"03ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"f0000000",
	x"00001fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffe00",
	x"03ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"f8000000",
	x"000003ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffe00",
	x"03ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"f8000000",
	x"00000000",
	x"00000fff",
	x"ffffffff",
	x"ffffffff",
	x"c0000000",
	x"00000000",
	x"00ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffe00",
	x"03ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fe000000",
	x"00000000",
	x"000000ff",
	x"ffffffff",
	x"ffffffff",
	x"00000000",
	x"00000000",
	x"000fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffe00",
	x"03ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ff000000",
	x"00000000",
	x"00000000",
	x"00000007",
	x"c0000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"03ffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffc00",
	x"03ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fff00000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"003fffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffc00",
	x"03ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffc0000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"0007ffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffc00",
	x"03ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"0001ffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffc00",
	x"03ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffff80",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000fff",
	x"ffffffff",
	x"ffffffff",
	x"fffffe00",
	x"03ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffe00000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000001",
	x"ffffffff",
	x"ffffffff",
	x"fffffe00",
	x"03ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fff80000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"7fffffff",
	x"ffffffff",
	x"fffffe00",
	x"03ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff8000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"3fffffff",
	x"ffffffff",
	x"fffffe00",
	x"03ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"1fffffff",
	x"ffffffff",
	x"fffffe00",
	x"03ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffff00",
	x"00180000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"00000000",
	x"1fffffff",
	x"ffffffff",
	x"fffffc00",
	x"03ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffe00",
	x"00000000",
	x"00000001",
	x"ffffffff",
	x"ffffffff",
	x"ffe00000",
	x"00000000",
	x"1fffffff",
	x"ffffffff",
	x"fffffc00",
	x"03ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffe0",
	x"00000000",
	x"0000000f",
	x"ffffffff",
	x"ffffffff",
	x"fffe0000",
	x"00000000",
	x"1fffffff",
	x"ffffffff",
	x"fffffc00",
	x"03ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"f8000000",
	x"1fffffff",
	x"ffffffff",
	x"fffff000",
	x"03ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fe000000",
	x"3fffffff",
	x"ffffffff",
	x"f8000000",
	x"03ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffc00000",
	x"7fffffff",
	x"ffffffff",
	x"e0000000",
	x"07ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffe00000",
	x"7fffffff",
	x"ffffffff",
	x"80000000",
	x"0fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffe00000",
	x"ffffffff",
	x"ffffffff",
	x"00000000",
	x"0fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffe00000",
	x"ffffffff",
	x"fffffffc",
	x"00000000",
	x"1fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffe00001",
	x"ffffffff",
	x"fffffff8",
	x"00000000",
	x"1fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffc00007",
	x"ffffffff",
	x"ffffffe0",
	x"00000000",
	x"3fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ff80000f",
	x"ffffffff",
	x"ffffff00",
	x"00000000",
	x"7fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fe00001f",
	x"ffffffff",
	x"fffff800",
	x"00000000",
	x"7fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fc00003f",
	x"ffffffff",
	x"ffff8000",
	x"00000000",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"f00000ff",
	x"ffffffff",
	x"fffc0000",
	x"00000001",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"e00001ff",
	x"ffffffff",
	x"fff00000",
	x"00000003",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"c00003ff",
	x"ffffffff",
	x"ff800000",
	x"00000007",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"80000fff",
	x"ffffffff",
	x"fe000000",
	x"0000000f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffffe",
	x"00001fff",
	x"ffffffff",
	x"f8000000",
	x"0000001f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffffc",
	x"00007fff",
	x"ffffffff",
	x"e0000000",
	x"0000007f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffff0",
	x"0000ffff",
	x"ffffffff",
	x"c0000000",
	x"7fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffe0",
	x"0001ffff",
	x"fffffff8",
	x"00000001",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffff00",
	x"0007ffff",
	x"ffffffc0",
	x"0000003f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffffc00",
	x"000fffff",
	x"fffff800",
	x"000001ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffff800",
	x"001fffff",
	x"fff80000",
	x"00000fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffe000",
	x"003fffff",
	x"fe000000",
	x"00007fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff8000",
	x"00ffffff",
	x"f0000000",
	x"0003ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffff0000",
	x"01ffffff",
	x"80000000",
	x"0007ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fffe0000",
	x"03fffffe",
	x"00000000",
	x"003fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fff80000",
	x"0ffffffc",
	x"00000000",
	x"00ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fff00000",
	x"1ffffff0",
	x"00000000",
	x"03ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffe00000",
	x"ffffffc0",
	x"00000000",
	x"07ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffc00003",
	x"ffffff80",
	x"00000000",
	x"3fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ff80000f",
	x"fffffe00",
	x"0000003f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ff00001f",
	x"fffffc00",
	x"000001ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ff00007f",
	x"fffff800",
	x"000fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fe0000ff",
	x"ffffe000",
	x"003fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"fc0000ff",
	x"ffffc000",
	x"00ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"f80001ff",
	x"ffff8000",
	x"01ffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"f00001ff",
	x"fffe0000",
	x"0fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"e00000ff",
	x"fff80000",
	x"3fffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"e00000ff",
	x"ffe00000",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"c000003f",
	x"fc000001",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"80000000",
	x"00000003",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"00000000",
	x"00000007",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"00000000",
	x"0000001f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"00000000",
	x"0000003f",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"00000000",
	x"000000ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"00000000",
	x"000001ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"00000000",
	x"000007ff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"80000000",
	x"00001fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"80000000",
	x"00007fff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"e0000000",
	x"0007ffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"f0000000",
	x"001fffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff",
	x"ffffffff"
	);	

begin
writing:	process(memwrite,clock)	
		begin	
		if(clock'event and clock='1')then
			if(MemWrite='1') then
			   RAM(conv_integer(address(31 downto 0)))<= write_data;
			end if;
		end if;
	end process;
read_data<=RAM(conv_integer(address(31 downto 0))) when memread='1' else x"00000000"; 
ext_read<=RAM(conv_integer(ext_addr(31 downto 0))); 
end  Behavioral;